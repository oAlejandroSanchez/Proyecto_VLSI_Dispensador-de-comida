--Arcvhivo que permite procesar la información del trigger

library ieee;
use ieee.std_logic_1164.all;

entity trigger is port(
	pwm,echo: in std_logic;
	salida: out std_logic);
end entity;

architecture arquitectura_trigger of trigger is
begin
	process(pwm)
	begin
		if(echo = '0') then
			salida <= pwm;
		end if;
	end process;
end architecture;